`include "modulos/nand.v"

module probadorTarea3 ();

initial begin
  $display("Modulo Probador de la Tarea 3");
end

endmodule
